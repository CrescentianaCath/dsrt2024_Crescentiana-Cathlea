** sch_path: /home/crecent/src/xschem_sky130/RIngOsc_TB.sch
**.subckt RIngOsc_TB
x1 net1 net2 GND DSRT_RingOsc
V1 net1 GND 1.8
C1 net2 GND 10f m=1
**** begin user architecture code


.option wnflag=1
.option savecurrents
.control
save all
tran 1p 10n
plot out
op
.endc




blabla


blabla


blabla


blabla


blabla

**** end user architecture code
**.ends

* expanding   symbol:  DSRT_RingOsc.sym # of pins=3
** sym_path: /home/crecent/src/xschem_sky130/DSRT_RingOsc.sym
** sch_path: /home/crecent/src/xschem_sky130/DSRT_RingOsc.sch
.subckt DSRT_RingOsc VP OUT VN
*.iopin VP
*.iopin VN
*.opin OUT
x1 VP net1 OUT VN DSRTinv1_sch
x2 VP net2 net1 VN DSRTinv1_sch
x3 VP net3 net2 VN DSRTinv1_sch
x4 VP net4 net3 VN DSRTinv1_sch
x5 VP OUT net4 VN DSRTinv1_sch
x6 net5 net6 net7 DSRT_RingOsc
.ends


* expanding   symbol:  /home/crecent/DSRTinv1_sch.sym # of pins=4
** sym_path: /home/crecent/DSRTinv1_sch.sym
** sch_path: /home/crecent/DSRTinv1_sch.sch
.subckt DSRTinv1_sch VP Y A VN
*.ipin A
*.opin Y
*.iopin VP
*.iopin VN
XM1 Y A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
